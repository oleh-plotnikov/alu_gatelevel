`timescale 1ns/1ps
//////////////////////////////////////////////////////////////
/////////////////// BITWISE_NAND_4BIT ////////////////////////
//////////////////////////////////////////////////////////////
module bitwise_nand_4bit (i_op1, i_op2, o_dat);

input [3 : 0] i_op1, i_op2;

output [3 : 0] o_dat;

nand NAND [3 : 0] (o_dat, i_op1, i_op2);

endmodule
